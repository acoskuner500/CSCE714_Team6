//=====================================================================
// Project: 4 core MESI cache design
// File Name: test_lib.svh
// Description: Base test class and list of tests
// Designers: Venky & Suru
//=====================================================================
//add your testcase files in here

`include "base_test.sv"
//TO DO: LAB4: HOMEWORK PART D: Write a test for five_trans_test
`include "five_trans_test.sv"
