//=====================================================================
// Project: 4 core MESI cache design
// File Name: test_lib.svh
// Description: Base test class and list of tests
// Designers: Venky & Suru
//=====================================================================
//add your testcase files in here

`include "base_test.sv"
`include "read_miss_icache.sv"
